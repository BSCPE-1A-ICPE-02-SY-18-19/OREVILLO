CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 8 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
76546066 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 49 296 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
317 0 0
2
5.89884e-315 0
0
2 +V
167 365 263 0 1 3
0 16
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3108 0 0
2
43530.4 0
0
2 +V
167 722 357 0 1 3
0 17
0
0 0 54256 180
3 10V
6 -2 27 6
3 V10
7 -12 28 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4299 0 0
2
43530.4 0
0
2 +V
167 537 357 0 1 3
0 18
0
0 0 54256 180
3 10V
6 -2 27 6
2 V9
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9672 0 0
2
43530.4 0
0
2 +V
167 366 358 0 1 3
0 19
0
0 0 54256 180
3 10V
6 -2 27 6
2 V8
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7876 0 0
2
43530.4 0
0
2 +V
167 216 356 0 1 3
0 20
0
0 0 54256 180
3 10V
6 -2 27 6
2 V7
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6369 0 0
2
43530.4 0
0
2 +V
167 722 261 0 1 3
0 21
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9172 0 0
2
43530.4 0
0
2 +V
167 537 261 0 1 3
0 22
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7100 0 0
2
43530.4 0
0
9 2-In AND~
219 630 136 0 3 22
0 15 12 14
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3820 0 0
2
43530.4 0
0
9 2-In AND~
219 441 127 0 3 22
0 10 11 15
0
0 0 624 0
5 74F08
-18 -24 17 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7678 0 0
2
43530.4 0
0
7 Pulser~
4 69 461 0 10 12
0 25 26 9 27 0 0 5 5 4
8
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
961 0 0
2
5.89884e-315 0
0
9 CC 7-Seg~
183 1092 71 0 18 19
10 8 7 5 6 4 3 2 9 28
0 0 1 1 1 1 1 1 2
0
0 0 21088 0
8 YELLOWCC
6 -41 62 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3178 0 0
2
5.89884e-315 0
0
6 74LS48
188 904 222 0 14 29
0 13 12 11 10 29 30 2 3 4
6 5 7 8 31
0
0 0 4848 0
6 74LS48
-21 -60 21 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3409 0 0
2
5.89884e-315 0
0
6 74112~
219 722 332 0 7 32
0 21 14 9 14 17 32 13
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 3 0
1 U
3951 0 0
2
5.89884e-315 0
0
6 74112~
219 537 332 0 7 32
0 22 15 9 15 18 33 12
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 3 0
1 U
8885 0 0
2
5.89884e-315 0
0
6 74112~
219 366 331 0 7 32
0 16 10 9 10 19 34 11
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
3780 0 0
2
5.89884e-315 0
0
6 74112~
219 215 331 0 7 32
0 23 24 9 24 20 35 10
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
9265 0 0
2
5.89884e-315 0
0
2 +V
167 216 261 0 1 3
0 23
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9442 0 0
2
5.89884e-315 0
0
36
7 7 2 0 0 8320 0 12 13 0 0 3
1107 107
1107 186
936 186
6 8 3 0 0 8320 0 12 13 0 0 3
1101 107
1101 195
936 195
5 9 4 0 0 8320 0 12 13 0 0 3
1095 107
1095 204
936 204
3 11 5 0 0 8320 0 12 13 0 0 3
1083 107
1083 222
936 222
4 10 6 0 0 8320 0 12 13 0 0 3
1089 107
1089 213
936 213
2 12 7 0 0 8320 0 12 13 0 0 3
1077 107
1077 231
936 231
1 13 8 0 0 8320 0 12 13 0 0 3
1071 107
1071 240
936 240
3 0 9 0 0 8192 0 17 0 0 12 3
185 304
162 304
162 452
3 0 9 0 0 0 0 16 0 0 12 3
336 304
324 304
324 452
3 0 9 0 0 0 0 15 0 0 12 3
507 305
487 305
487 452
3 0 9 0 0 0 0 14 0 0 12 3
692 305
677 305
677 452
3 8 9 0 0 4224 0 11 12 0 0 3
93 452
1113 452
1113 107
4 0 10 0 0 12416 0 13 0 0 34 5
872 213
802 213
802 396
254 396
254 295
3 0 11 0 0 12416 0 13 0 0 23 5
872 204
793 204
793 387
407 387
407 294
2 0 12 0 0 12416 0 13 0 0 19 5
872 195
782 195
782 377
574 377
574 294
1 7 13 0 0 8320 0 13 14 0 0 4
872 186
773 186
773 296
746 296
2 0 14 0 0 4096 0 14 0 0 18 2
698 296
665 296
3 4 14 0 0 8320 0 9 14 0 0 4
651 136
665 136
665 314
698 314
2 7 12 0 0 0 0 9 15 0 0 4
606 145
574 145
574 296
561 296
2 0 15 0 0 4096 0 15 0 0 21 2
513 296
477 296
4 0 15 0 0 8320 0 15 0 0 22 3
513 314
477 314
477 127
3 1 15 0 0 0 0 10 9 0 0 2
462 127
606 127
2 7 11 0 0 0 0 10 16 0 0 4
417 136
407 136
407 295
390 295
1 0 10 0 0 0 0 10 0 0 33 3
417 118
312 118
312 296
1 1 16 0 0 4224 0 2 16 0 0 3
365 272
365 268
366 268
1 5 17 0 0 4224 0 3 14 0 0 2
722 342
722 344
1 5 18 0 0 4224 0 4 15 0 0 2
537 342
537 344
1 5 19 0 0 0 0 5 16 0 0 2
366 343
366 343
1 5 20 0 0 4224 0 6 17 0 0 3
216 341
216 343
215 343
1 1 21 0 0 4224 0 7 14 0 0 2
722 270
722 269
1 1 22 0 0 4224 0 8 15 0 0 2
537 270
537 269
1 1 23 0 0 4224 0 18 17 0 0 3
216 270
216 268
215 268
4 0 10 0 0 0 0 16 0 0 34 3
342 313
312 313
312 295
7 2 10 0 0 0 0 17 16 0 0 2
239 295
342 295
4 0 24 0 0 4096 0 17 0 0 36 3
191 313
118 313
118 295
1 2 24 0 0 8320 0 1 17 0 0 3
61 296
61 295
191 295
2
-24 0 0 0 400 255 0 0 0 3 2 1 66
13 Comic Sans MS
0 0 0 26
12 558 424 610
28 567 407 603
26 EUNEROSE OREVILLO BSCpE 1A
-24 0 0 0 400 255 0 0 0 3 2 1 18
8 Elephant
0 0 0 25
68 28 565 75
84 37 548 68
25 4-BIT SYNCHRONOUS COUNTER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
